library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use ieee.math_real.ceil;
    use ieee.math_real.floor;
    use ieee.math_real.log2;
    use std.env.finish;
    use std.env.stop;
    use std.textio.all;

library accel;
    use accel.utilities.all;

entity kernels_tb is
    generic (
        size_x : positive := 7;
        size_y : positive := 10;

        line_length_iact : positive := 32; /* TODO check influence on tiling - does not work for length 32, kernel 4 and channels 10. Does not work for length 30, kernel 3 and channels 10*/
        line_length_psum : positive := 128;
        line_length_wght : positive := 32; /* TODO check influence on tiling - does not work for length 32, kernel 4 and channels 10. Does not work for length 30, kernel 3 and channels 10*/

        data_width_input : positive := 8;  -- Width of the input data (weights, iacts)
        data_width_psum  : positive := 16; -- or 17??

        mem_word_count : positive := 8;
        mem_addr_width : positive := 15;

        g_channels    : positive := 8;
        g_image_y     : positive := 16;
        g_image_x     : positive := 16;
        g_kernel_size : positive := 5;

        g_iact_fifo_size : positive := 15;
        g_wght_fifo_size : positive := 15;
        g_psum_fifo_size : positive := 128;

        g_clk    : time := 10000 ps; -- ps
        g_clk_sp : time := 1000 ps;  -- ps

        g_files_dir : string  := "test/image_size_16_kernel_size_5_c_8/";
        g_init_sp   : boolean := true;

        -- g_h2 : positive := positive(integer(ceil(real(g_image_x - g_kernel_size + 1) / real(size_x)))); -- Y tiles, determined in control module, but for input data loading required here
        g_h2 : positive := positive(integer(ceil(real(g_image_x) / real(size_x)))); -- Y tiles, determined in control module, but for input data loading required here
        g_m0 : positive := positive(integer(floor(real(size_y) / real(g_kernel_size))))
    );
end entity kernels_tb;

architecture imp of kernels_tb is

    constant size_rows      : positive := size_x + size_y - 1;
    constant mem_data_width : positive := mem_word_count * data_width_input;

    signal clk    : std_logic := '0';
    signal clk_sp : std_logic := '0';
    signal rstn   : std_logic;

    signal start, done : std_logic;

    signal o_psums           : array_t(0 to size_x - 1)(data_width_psum - 1 downto 0);
    signal o_psums_valid     : std_logic_vector(size_x - 1 downto 0);
    signal i_data_iact       : array_t (0 to size_rows - 1)(data_width_input - 1 downto 0);
    signal i_data_iact_valid : std_logic_vector(size_rows - 1 downto 0);
    signal i_data_wght       : array_t (0 to size_y - 1)(data_width_input - 1 downto 0);
    signal i_data_wght_valid : std_logic_vector(size_y - 1 downto 0);

    signal s_input_image     : int_image_t(0 to size_rows - 1, 0 to g_image_x * g_channels * g_h2 - 1);         -- 2, because two tile_y
    signal s_input_weights   : int_image_t(0 to g_kernel_size - 1, 0 to g_kernel_size * g_channels * g_h2 - 1); -- not *2 because kernel stays the same across tile_y
    signal s_expected_output : int_image_t(0 to g_image_y - g_kernel_size, 0 to g_image_x - g_kernel_size);

    signal write_en_iact : std_logic;
    signal write_en_wght : std_logic;
    signal din_iact      : std_logic_vector(data_width_input - 1 downto 0);
    signal din_wght      : std_logic_vector(data_width_input - 1 downto 0);

    signal w_h2 : integer;
    signal w_m0 : integer;

    type   ram_type is array (0 to 2 ** mem_addr_width / mem_word_count - 1) of std_logic_vector(mem_data_width - 1 downto 0);
    type   ram_cols_type is array(0 to mem_word_count) of ram_type;
    signal ram_cols : ram_cols_type;

    type t_state is (s_calculate, s_output, s_incr_c1);

    signal params : parameters_t := (
                                     kernel_size => g_kernel_size,
                                     image_x => g_image_x,
                                     image_y => g_image_y,
                                     inputchs => g_channels,
                                     w1 => g_image_x,
                                     m0 => 1,
                                     requant_enab => false,
                                     mode_act => passthrough,
                                     mode_pad => none,
                                     bias => (others => 0),
                                     zeropt_fp32 => (others => (others => '0')),
                                     scale_fp32 => (others => (others => '0')),
                                     others => 0
                                    );

begin

    o_psums           <= << signal accelerator_inst.w_psums : array_t(0 to size_x - 1)(data_width_psum - 1 downto 0) >>;
    o_psums_valid     <= << signal accelerator_inst.w_psums_valid : std_logic_vector(size_x - 1 downto 0) >>;
    i_data_iact       <= << signal accelerator_inst.w_data_iact : array_t (0 to size_rows - 1)(data_width_input - 1 downto 0) >>;
    i_data_iact_valid <= << signal accelerator_inst.w_data_iact_valid : std_logic_vector(size_rows - 1 downto 0) >>;
    i_data_wght       <= << signal accelerator_inst.w_data_wght : array_t (0 to size_y - 1)(data_width_input - 1 downto 0) >>;
    i_data_wght_valid <= << signal accelerator_inst.w_data_wght_valid : std_logic_vector(size_y - 1 downto 0) >>;

    w_h2 <= << signal accelerator_inst.w_h2 : integer >>;
    w_m0 <= << signal accelerator_inst.w_m0 : integer >>;

    write_en_iact <= '0';
    write_en_wght <= '0';
    din_iact      <= (others => '0');
    din_wght      <= (others => '0');

    accelerator_inst : entity work.accelerator
        generic map (
            size_x           => size_x,
            size_y           => size_y,
            line_length_iact => line_length_iact,
            line_length_wght => line_length_wght,
            line_length_psum => line_length_psum,
            data_width_input => data_width_input,
            data_width_psum  => data_width_psum
        )
        port map (
            clk            => clk,
            rstn           => rstn,
            clk_sp         => clk_sp,
            i_start        => start,
            o_done         => done,
            i_params       => params,
            o_status       => open,
            i_mem_en       => '0',
            i_mem_write_en => (others => '0'),
            i_mem_addr     => (others => '0'),
            i_mem_din      => (others => '0')
        );

    rstn_gen : process is
    begin

        rstn  <= '0';
        start <= '0';
        wait for 100 ns;
        rstn  <= '1';
        wait for 20 ns;
        start <= '1';
        wait;

    end process rstn_gen;

    clk_gen : process (clk) is
    begin

        clk <= not clk after g_clk;

    end process clk_gen;

    clk_sp_gen : process (clk_sp) is
    begin

        clk_sp <= not clk_sp after g_clk_sp;

    end process clk_sp_gen;

    p_constant_check : process is
    begin

        -- assert line_length_iact >= g_kernel_size * g_channels
        --     report "Line length to store input values must be greater or equal to the kernel size"
        --     severity failure;

        assert size_y >= g_kernel_size
            report "Y dimension of PE array has to be greater or equal to kernel size"
            severity failure;

        -- assert line_length_wght >= g_kernel_size * g_channels
        --     report "Length of wght buffer has to be greater or equal to kernel size, buffer has to store values of one kernel row at a time."
        --     severity failure;

        assert line_length_psum >= g_image_x - g_kernel_size
            report "Psum buffer has to hold output values of one row, must not be smaller than output row size"
            severity failure; /* TODO To be changed by splitting the task and propagating as many psums that the buffer can hold through the array at once */

        wait;

    end process p_constant_check;

    p_read_files : process is
    begin

        s_input_image <= read_file(file_name => g_files_dir & "_image_reordered_2.txt", num_col => g_image_x * g_channels * g_h2, num_row => size_rows);
        -- s_input_weights   <= read_file(file_name => "src/_kernel_reordered.txt", num_col => g_kernel_size * g_channels * g_tiles_y, num_row => g_kernel_size);
        s_expected_output <= read_file(file_name => g_files_dir & "_convolution.txt", num_col => g_image_x - g_kernel_size + 1, num_row => g_image_y - g_kernel_size + 1);
        wait;

    end process p_read_files;

    p_check_img : for y in 0 to size_rows - 1 generate

        p_check_image_vals : process is
        begin

            for i in 0 to g_image_x * g_channels * g_h2 - 1 loop

                wait until rising_edge(clk) and i_data_iact_valid(y) = '1';

                if i_data_iact(y) /= std_logic_vector(to_signed(s_input_image(y, i), data_width_input)) then
                    assert i_data_iact(y) = std_logic_vector(to_signed(s_input_image(y, i), data_width_input))
                        report "Input iact " & integer'image(i) & " wrong. Iact is " & integer'image(to_integer(signed(i_data_iact(y)))) & " - should be "
                               & integer'image(s_input_image(y, i))
                        severity warning;
                else
                -- report "Got correct iact " & integer'image(to_integer(signed(i_data_iact(y)))) & " (" & integer'image(i) & ")";
                end if;

            end loop;

            while true loop

                assert i_data_iact_valid(y) = '0'
                    report "Input data iact should not be valid!"
                    severity warning;

                wait until i_data_iact_valid(y)'event;

            end loop;

        end process p_check_image_vals;

    end generate p_check_img;

    /*p_check_wght : for y in 0 to size_y - 1 generate

        p_check_wght_vals : process is
        begin

            for i in 0 to g_kernel_size * g_channels * g_tiles_y - 1 loop

                wait until rising_edge(clk) and i_data_wght_valid(y) = '1';

                assert i_data_wght(y) = std_logic_vector(to_signed(s_input_weights(y, i), data_width_input))
                    report "Input wght (" & integer'image(y) & ") wrong. Wght is " & integer'image(to_integer(signed(i_data_wght(y)))) & " - should be "
                           & integer'image(s_input_weights(y, i))
                    severity warning;

                report "Got correct (" & integer'image(y) & ") wght " & integer'image(to_integer(signed(i_data_wght(y))));

            end loop;

            while true loop

                assert i_data_wght_valid(y) = '0'
                    report "Input data wght should not be valid!"
                    severity warning;

                wait until i_data_wght_valid(y)'event;

            end loop;

        end process p_check_wght_vals;

    end generate p_check_wght;*/

    write_outputs : process is

        file     outfile : text open write_mode is g_files_dir & "_output.txt";
        variable row     : line;

    begin

        wait until done = '1';

        wait for 2000 ns;

        -- TODO: fix writeout for multi-column spad
        for i in 0 to 2 ** mem_addr_width / mem_word_count - 1 loop

            write(row, integer'image(to_integer(signed(ram_cols(0)(i)))));
            writeline(outfile, row);

        end loop;

        report "Writing outputs is finished."
            severity note;
        finish;

        wait;

    end process write_outputs;

    -- assemble all scratchpad columns into ram_cols for easy access

    gen_ram_alias : for i in 0 to mem_word_count - 1 generate

        ram_alias : process is

            alias ram is << variable ^.accelerator_inst.scratchpad_inst.ram.gen_cols(i).ram.ram : ram_type >>;

        begin

            wait until done = '1';
            wait for 900 ns;
            ram_cols(i) <= ram;
            wait;

        end process ram_alias;

    end generate gen_ram_alias;

end architecture imp;
