library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;
    use work.utilities.all;

entity pe_array is
    generic (

    );
    port (
        clk  : in    std_logic;
        rstn : in    std_logic;


    );
end entity pe_array;

architecture behavioral of pe_array is
begin

end architecture behavioral;